../../integration/tb/bootrom_64.sv