module culsans_tb ();

// Clock generator

// Reset generator

// Detect the end of the simulation

// DUT

// ...

endmodule
