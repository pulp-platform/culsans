module xlnx_ila(clk, probe0, probe1, probe2, probe3, probe4, probe5, 
                probe6, probe7, probe8, probe9, probe10, probe11, probe12);
   
  input clk;
   input [31:0] probe0;
   input [31:0] probe1;
   input [31:0] probe2;
   input [31:0] probe3;
   input [31:0] probe4;
   input [31:0] probe5;
   input [31:0] probe6;
   input [31:0] probe7;
   input [31:0] probe8;
   input [31:0] probe9;
   input [31:0] probe10;
   input [31:0] probe11;
   input [47:0] probe12;
endmodule
