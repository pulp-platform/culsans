../../integration/tb/ila.sv